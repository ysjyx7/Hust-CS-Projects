/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : ROM_ROM                                                      **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module ROM_ROM( Address,
                Data);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input[9:0]  Address;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] Data;
   reg[31:0] Data;

   always @ (Address)
   begin
      case(Address)
0 : Data = 32'h03000713;
1 : Data = 32'h00000593;
2 : Data = 32'h02200513;
3 : Data = 32'h00000073;
4 : Data = 32'h02300513;
5 : Data = 32'h00000073;
6 : Data = 32'h02060063;
7 : Data = 32'h40e60633;
8 : Data = 32'h00058793;
9 : Data = 32'h00359593;
10 : Data = 32'h00f585b3;
11 : Data = 32'h00f585b3;
12 : Data = 32'h00c585b3;
13 : Data = 32'hfc000ee3;
14 : Data = 32'h00000693;
15 : Data = 32'h02200513;
16 : Data = 32'h00000073;
17 : Data = 32'h02300513;
18 : Data = 32'h00000073;
19 : Data = 32'h02060063;
20 : Data = 32'h40e60633;
21 : Data = 32'h00068793;
22 : Data = 32'h00369693;
23 : Data = 32'h00f686b3;
24 : Data = 32'h00f686b3;
25 : Data = 32'h00c686b3;
26 : Data = 32'hfc000ee3;
27 : Data = 32'h02b68663;
28 : Data = 32'h00b6ec63;
29 : Data = 32'h00000263;
30 : Data = 32'h00d00513;
31 : Data = 32'h0db00893;
32 : Data = 32'h00000073;
33 : Data = 32'hfa000ae3;
34 : Data = 32'h00d00513;
35 : Data = 32'h03200893;
36 : Data = 32'h00000073;
37 : Data = 32'hfa0002e3;
38 : Data = 32'h00d00513;
39 : Data = 32'h03600893;
40 : Data = 32'h00000073;
41 : Data = 32'hf60000e3;


         default : Data = 0;
      endcase
   end

endmodule
