/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : Bit_Extender_2_5_SIGN                                        **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module Bit_Extender_2_5_SIGN( imm_in,
                              imm_out);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input[1:0]  imm_in;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output reg [4:0] imm_out;

	always @(*) begin
		imm_out = {{(3){imm_in[1]}}, imm_in};
	end

endmodule
