/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : LogisimCounter                                               **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module LogisimCounter(clk,enable,Q);

   /***************************************************************************
    ** Here all module parameters are defined with a dummy value             **
    ***************************************************************************/
  

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input clk,enable;
   output [31:0]Q;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   reg [31:0]cnt;
   initial
   begin
   cnt=0;
   end
assign Q=cnt;
   /***************************************************************************
    ** Functionality of the counter:                                         **
    ** __Load_Count_|_mode                                                   **
    ** ____0____0___|_halt                                                   **
    ** ____0____1___|_count_up_(default)                                     **
    ** ____1____0___|load                                                    **
    ** ____1____1___|_count_down                                             **
    ***************************************************************************/

 always @(posedge clk)
begin
   if(enable)
   begin
   cnt<=cnt+1;
   end
end



endmodule
